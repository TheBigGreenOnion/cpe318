library ieee;
use ieee.std_logic_1164.all;

entity  is
    port ( ); 
end entity ;

architecture verify of  is
    signal 
begin
    duv : entity work.
        port map ( );

    test : process is
    begin

end architecture verify;
